// File:    kernel_sum.sv
// Author:  Lei Kuang
// Date:    20th of August 2019
// @ Imperial College London

module kernel_sum_tb;

logic        clk;
logic [31:0] kernel [48:0];
logic        kernel_valid;
logic [31:0] sum;
logic        sum_valid;

kernel_sum kernel_sum_inst(.*);

initial begin
    clk = '0;
    forever #2.5ns clk = ~clk;
end

initial begin
    kernel_valid = '0;
    
    @(posedge clk)
    #1ns kernel_valid = '1;
    @(posedge clk)
    #1ns kernel_valid = '0;
    
    @(posedge clk)
    #1ns kernel_valid = '1;
    @(posedge clk)
    #1ns kernel_valid = '0;
    
    @(posedge clk)
    #1ns kernel_valid = '1;
    @(posedge clk)
    #1ns kernel_valid = '1;
    @(posedge clk)
    #1ns kernel_valid = '0;
end

assign kernel [ 0] = 32'b00111011100101001110010011011101;
assign kernel [ 1] = 32'b00111011111111110110110001011101;
assign kernel [ 2] = 32'b00111100010000111101010111100011;
assign kernel [ 3] = 32'b00111100011100100011001111100100;
assign kernel [ 4] = 32'b00111100000111110011000000110010;
assign kernel [ 5] = 32'b00111100000011011011011110111111;
assign kernel [ 6] = 32'b00111011100101111011011001001100;
assign kernel [ 7] = 32'b00111100000101011110101011111000;
assign kernel [ 8] = 32'b00111100001011101111111110000010;
assign kernel [ 9] = 32'b00111100101001011100100011100101;
assign kernel [10] = 32'b00111100111010000000110000001110;
assign kernel [11] = 32'b00111100101000000100100001101011;
assign kernel [12] = 32'b00111100011101010011111111001111;
assign kernel [13] = 32'b00111011111011111111001010101111;
assign kernel [14] = 32'b00111100010110101001101101011011;
assign kernel [15] = 32'b00111100110011000011010010101000;
assign kernel [16] = 32'b00111100110101000000001001000001;
assign kernel [17] = 32'b00111101000110100011110001001001;
assign kernel [18] = 32'b00111101000000000001000011001111;
assign kernel [19] = 32'b00111100101101101110111100110111;
assign kernel [20] = 32'b00111100010110110011100011111010;
assign kernel [21] = 32'b00111011110001111011101111001111;
assign kernel [22] = 32'b00111100101010111101100111011011;
assign kernel [23] = 32'b00111101000110100011110001001001;
assign kernel [24] = 32'b00111101001111110100101001011101;
assign kernel [25] = 32'b00111101001010000101011011010001;
assign kernel [26] = 32'b00111100001101000101001111011011;
assign kernel [27] = 32'b00111100001110111000001011010000;
assign kernel [28] = 32'b00111011111111001010010100010100;
assign kernel [29] = 32'b00111100100101111010100001110001;
assign kernel [30] = 32'b00111100110010110010111111101101;
assign kernel [31] = 32'b00111101001001010111100001110101;
assign kernel [32] = 32'b00111101000101001100101010000100;
assign kernel [33] = 32'b00111100110011001000011001101000;
assign kernel [34] = 32'b00111100001010001000111010100011;
assign kernel [35] = 32'b00111011111100111111010010001000;
assign kernel [36] = 32'b00111100100010111010010111111101;
assign kernel [37] = 32'b00111100101101101110111100110111;
assign kernel [38] = 32'b00111100110101000000001001000001;
assign kernel [39] = 32'b00111100101111101110000001110001;
assign kernel [40] = 32'b00111100100000001001011100000000;
assign kernel [41] = 32'b00111011111010111101101111101111;
assign kernel [42] = 32'b00111011100101111011011001001100;
assign kernel [43] = 32'b00111011101011011010001111011101;
assign kernel [44] = 32'b00111100010101011011111000111110;
assign kernel [45] = 32'b00111100011110000101010110000111;
assign kernel [46] = 32'b00111100010110100010000100010010;
assign kernel [47] = 32'b00111100000101101001111101001011;
assign kernel [48] = 32'b00111011011001011000100111000101;

endmodule
