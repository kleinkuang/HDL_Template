// File:    kernel_product_tb.sv
// Author:  Lei Kuang
// Date:    21th of August 2019
// @ Imperial College London

module kernel_product_tb;

logic        clk                ;
logic [31:0] kernel_a [48:0]    ;
logic [31:0] kernel_b [48:0]    ;
logic        kernel_valid       ;
logic [31:0] product [48:0]     ;
logic        product_valid      ;

kernel_product kernel_product_inst(.*);

initial begin
    clk = '0;
    forever #2.5ns clk = ~clk;
end

initial begin
    kernel_valid = '0;
    @(posedge clk)
    for(int i=0; i<5; i++) begin
        @(negedge clk)
        kernel_valid = '1;
        @(negedge clk)
        kernel_valid = '0;
    end
end

assign kernel_a [ 0] = 32'b00111011101000010100101110000010;
assign kernel_a [ 1] = 32'b00111100000101101010101101011001;
assign kernel_a [ 2] = 32'b00111100010110110011100011111011;
assign kernel_a [ 3] = 32'b00111100011110000110100101100110;
assign kernel_a [ 4] = 32'b00111100010110110011100011111011;
assign kernel_a [ 5] = 32'b00111100000101101010101101011001;
assign kernel_a [ 6] = 32'b00111011101000010100101110000010;
assign kernel_a [ 7] = 32'b00111100000101101010101101011001;
assign kernel_a [ 8] = 32'b00111100100011001011111001100010;
assign kernel_a [ 9] = 32'b00111100110011001100011111100110;
assign kernel_a [10] = 32'b00111100111010000000110000001110;
assign kernel_a [11] = 32'b00111100110011001100011111100110;
assign kernel_a [12] = 32'b00111100100011001011111001100010;
assign kernel_a [13] = 32'b00111100000101101010101101011001;
assign kernel_a [14] = 32'b00111100010110110011100011111011;
assign kernel_a [15] = 32'b00111100110011001100011111100110;
assign kernel_a [16] = 32'b00111101000101001111101000101001;
assign kernel_a [17] = 32'b00111101001010001101000000110010;
assign kernel_a [18] = 32'b00111101000101001111101000101001;
assign kernel_a [19] = 32'b00111100110011001100011111100110;
assign kernel_a [20] = 32'b00111100010110110011100011111011;
assign kernel_a [21] = 32'b00111100011110000110100101100110;
assign kernel_a [22] = 32'b00111100111010000000110000001110;
assign kernel_a [23] = 32'b00111101001010001101000000110010;
assign kernel_a [24] = 32'b00111101001111110100101001011101;
assign kernel_a [25] = 32'b00111101001010001101000000110010;
assign kernel_a [26] = 32'b00111100111010000000110000001110;
assign kernel_a [27] = 32'b00111100011110000110100101100110;
assign kernel_a [28] = 32'b00111100010110110011100011111011;
assign kernel_a [29] = 32'b00111100110011001100011111100110;
assign kernel_a [30] = 32'b00111101000101001111101000101001;
assign kernel_a [31] = 32'b00111101001010001101000000110010;
assign kernel_a [32] = 32'b00111101000101001111101000101001;
assign kernel_a [33] = 32'b00111100110011001100011111100110;
assign kernel_a [34] = 32'b00111100010110110011100011111011;
assign kernel_a [35] = 32'b00111100000101101010101101011001;
assign kernel_a [36] = 32'b00111100100011001011111001100010;
assign kernel_a [37] = 32'b00111100110011001100011111100110;
assign kernel_a [38] = 32'b00111100111010000000110000001110;
assign kernel_a [39] = 32'b00111100110011001100011111100110;
assign kernel_a [40] = 32'b00111100100011001011111001100010;
assign kernel_a [41] = 32'b00111100000101101010101101011001;
assign kernel_a [42] = 32'b00111011101000010100101110000010;
assign kernel_a [43] = 32'b00111100000101101010101101011001;
assign kernel_a [44] = 32'b00111100010110110011100011111011;
assign kernel_a [45] = 32'b00111100011110000110100101100110;
assign kernel_a [46] = 32'b00111100010110110011100011111011;
assign kernel_a [47] = 32'b00111100000101101010101101011001;
assign kernel_a [48] = 32'b00111011101000010100101110000010;

assign kernel_b [ 0] = 32'b00111111010100101001010001110010;
assign kernel_b [ 1] = 32'b00111111010101011101010001000101;
assign kernel_b [ 2] = 32'b00111110110000000010100011000110;
assign kernel_b [ 3] = 32'b00111110110000000010100011000110;
assign kernel_b [ 4] = 32'b00111111010101011101010001000101;
assign kernel_b [ 5] = 32'b00111111010100101001010001110010;
assign kernel_b [ 6] = 32'b00111111011111111110101110000110;
assign kernel_b [ 7] = 32'b00111110110011011101010110111111;
assign kernel_b [ 8] = 32'b00111110110110111110111011110001;
assign kernel_b [ 9] = 32'b00111111011000011110101101010001;
assign kernel_b [10] = 32'b00111111011000011110101101010001;
assign kernel_b [11] = 32'b00111110110110111110111011110001;
assign kernel_b [12] = 32'b00111110110011011101010110111111;
assign kernel_b [13] = 32'b00111111011011000101000101011010;
assign kernel_b [14] = 32'b00111111010100101001010001110010;
assign kernel_b [15] = 32'b00111111011111111110101110000110;
assign kernel_b [16] = 32'b00111111100000000000000000000000;
assign kernel_b [17] = 32'b00111111100000000000000000000000;
assign kernel_b [18] = 32'b00111111011111111110101110000110;
assign kernel_b [19] = 32'b00111111010100101001010001110010;
assign kernel_b [20] = 32'b00111111001101100010100000000001;
assign kernel_b [21] = 32'b00111111010100101001010001110010;
assign kernel_b [22] = 32'b00111111011111111110101110000110;
assign kernel_b [23] = 32'b00111111100000000000000000000000;
assign kernel_b [24] = 32'b00111111100000000000000000000000;
assign kernel_b [25] = 32'b00111111011111111110101110000110;
assign kernel_b [26] = 32'b00111111010100101001010001110010;
assign kernel_b [27] = 32'b00111111001101100010100000000001;
assign kernel_b [28] = 32'b00111110110011011101010110111111;
assign kernel_b [29] = 32'b00111110110110111110111011110001;
assign kernel_b [30] = 32'b00111111011000011110101101010001;
assign kernel_b [31] = 32'b00111111011000011110101101010001;
assign kernel_b [32] = 32'b00111110110110111110111011110001;
assign kernel_b [33] = 32'b00111110110011011101010110111111;
assign kernel_b [34] = 32'b00111111011011000101000101011010;
assign kernel_b [35] = 32'b00111111010100101001010001110010;
assign kernel_b [36] = 32'b00111111010101011101010001000101;
assign kernel_b [37] = 32'b00111110110000000010100011000110;
assign kernel_b [38] = 32'b00111110110000000010100011000110;
assign kernel_b [39] = 32'b00111111010101011101010001000101;
assign kernel_b [40] = 32'b00111111010100101001010001110010;
assign kernel_b [41] = 32'b00111111011111111110101110000110;
assign kernel_b [42] = 32'b00111111011110000001111110101011;
assign kernel_b [43] = 32'b00111111001110011110010011101000;
assign kernel_b [44] = 32'b00111111100000000000000000000000;
assign kernel_b [45] = 32'b00111111100000000000000000000000;
assign kernel_b [46] = 32'b00111111001110011110010011101000;
assign kernel_b [47] = 32'b00111111011110000001111110101011;
assign kernel_b [48] = 32'b00111111011111110100011111110000;

endmodule
