// File:    gaussian_kernel.sv
// Author:  Lei Kuang
// Date:    20th of August 2019
// @ Imperial College London

module gaussian_kernel
(
    output logic [31:0] gaussian_kernel [48:0]
);

// By Matlab
/*
% Pre-compute space weights (unchanged)
[x,y] = meshgrid(-r:r,-r:r);
D = exp(-(x.^2+y.^2)/(2*sigma_s^2));
% Normalization
D = D ./ sum(D(:));
% Gaussian Kernel
for i=1:7
    for j=1:7
        fprintf('assign weights [%2d] = 64''b%s;\n', i*7+j-8, dec2bin(typecast(D(i,j), 'uint64'),64));
    end
end
*/

assign gaussian_kernel [ 0] = 32'b00111011101000010100101110000010;
assign gaussian_kernel [ 1] = 32'b00111100000101101010101101011001;
assign gaussian_kernel [ 2] = 32'b00111100010110110011100011111011;
assign gaussian_kernel [ 3] = 32'b00111100011110000110100101100110;
assign gaussian_kernel [ 4] = 32'b00111100010110110011100011111011;
assign gaussian_kernel [ 5] = 32'b00111100000101101010101101011001;
assign gaussian_kernel [ 6] = 32'b00111011101000010100101110000010;
assign gaussian_kernel [ 7] = 32'b00111100000101101010101101011001;
assign gaussian_kernel [ 8] = 32'b00111100100011001011111001100010;
assign gaussian_kernel [ 9] = 32'b00111100110011001100011111100110;
assign gaussian_kernel [10] = 32'b00111100111010000000110000001110;
assign gaussian_kernel [11] = 32'b00111100110011001100011111100110;
assign gaussian_kernel [12] = 32'b00111100100011001011111001100010;
assign gaussian_kernel [13] = 32'b00111100000101101010101101011001;
assign gaussian_kernel [14] = 32'b00111100010110110011100011111011;
assign gaussian_kernel [15] = 32'b00111100110011001100011111100110;
assign gaussian_kernel [16] = 32'b00111101000101001111101000101001;
assign gaussian_kernel [17] = 32'b00111101001010001101000000110010;
assign gaussian_kernel [18] = 32'b00111101000101001111101000101001;
assign gaussian_kernel [19] = 32'b00111100110011001100011111100110;
assign gaussian_kernel [20] = 32'b00111100010110110011100011111011;
assign gaussian_kernel [21] = 32'b00111100011110000110100101100110;
assign gaussian_kernel [22] = 32'b00111100111010000000110000001110;
assign gaussian_kernel [23] = 32'b00111101001010001101000000110010;
assign gaussian_kernel [24] = 32'b00111101001111110100101001011101;
assign gaussian_kernel [25] = 32'b00111101001010001101000000110010;
assign gaussian_kernel [26] = 32'b00111100111010000000110000001110;
assign gaussian_kernel [27] = 32'b00111100011110000110100101100110;
assign gaussian_kernel [28] = 32'b00111100010110110011100011111011;
assign gaussian_kernel [29] = 32'b00111100110011001100011111100110;
assign gaussian_kernel [30] = 32'b00111101000101001111101000101001;
assign gaussian_kernel [31] = 32'b00111101001010001101000000110010;
assign gaussian_kernel [32] = 32'b00111101000101001111101000101001;
assign gaussian_kernel [33] = 32'b00111100110011001100011111100110;
assign gaussian_kernel [34] = 32'b00111100010110110011100011111011;
assign gaussian_kernel [35] = 32'b00111100000101101010101101011001;
assign gaussian_kernel [36] = 32'b00111100100011001011111001100010;
assign gaussian_kernel [37] = 32'b00111100110011001100011111100110;
assign gaussian_kernel [38] = 32'b00111100111010000000110000001110;
assign gaussian_kernel [39] = 32'b00111100110011001100011111100110;
assign gaussian_kernel [40] = 32'b00111100100011001011111001100010;
assign gaussian_kernel [41] = 32'b00111100000101101010101101011001;
assign gaussian_kernel [42] = 32'b00111011101000010100101110000010;
assign gaussian_kernel [43] = 32'b00111100000101101010101101011001;
assign gaussian_kernel [44] = 32'b00111100010110110011100011111011;
assign gaussian_kernel [45] = 32'b00111100011110000110100101100110;
assign gaussian_kernel [46] = 32'b00111100010110110011100011111011;
assign gaussian_kernel [47] = 32'b00111100000101101010101101011001;
assign gaussian_kernel [48] = 32'b00111011101000010100101110000010;

endmodule
